{%- import "utils_tmpl.sv" as utils with context -%}


{{hwif.get_package_declaration()}}

