{%- filter indent %}
{%- block body %}
{%- endblock %}
{%- endfilter %}
